LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;

ENTITY VGA_CONTROLLER IS
	PORT(
		SW : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		KEY : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
		CLOCK_50 : IN STD_LOGIC;
		LEDG : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		DRAM_CLK, DRAM_CKE : OUT STD_LOGIC;
		DRAM_ADDR : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
		DRAM_BA_0, DRAM_BA_1 : BUFFER STD_LOGIC;
		DRAM_CS_N, DRAM_CAS_N, DRAM_RAS_N, DRAM_WE_N : OUT STD_LOGIC;
		DRAM_DQ : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		DRAM_UDQM, DRAM_LDQM : BUFFER STD_LOGIC;
		
		VGA_R:out	std_logic_vector(9	downto	0);	
		VGA_G:out	std_logic_vector(9	downto	0);	
		VGA_B:out	std_logic_vector(9	downto	0);	
		VGA_CLK:	out	std_logic;
		VGA_BLANK:	out	std_logic;	
		VGA_HS:out	std_logic;	
		VGA_VS:out	std_logic;	
		VGA_SYNC:out	std_logic;
		SRAM_DQ	:	INOUT	STD_LOGIC_VECTOR(15	downto	0);
		SRAM_ADDR	:	OUT	STD_LOGIC_VECTOR(17	downto	0);
		SRAM_LB_N	:	OUT	STD_LOGIC;
		SRAM_UB_N	:	OUT	STD_LOGIC;
		SRAM_CE_N	:	OUT	STD_LOGIC;
		SRAM_OE_N	:	OUT	STD_LOGIC;
		SRAM_WE_N	:	OUT	STD_LOGIC
	);
END VGA_CONTROLLER;

ARCHITECTURE STRUCTURE OF VGA_CONTROLLER IS
component VGA_GRAPHICS is
        port (
            clk_clk                                         : in    std_logic;                     		  	          -- clk
            reset_reset_n                                   : in    std_logic;                                        -- reset_n
            sdram_wire_addr                                 : out   std_logic_vector(11 downto 0);                    -- addr
            sdram_wire_ba                                   : out   std_logic_vector(1 downto 0);                     -- ba
            sdram_wire_cas_n                                : out   std_logic;                                        -- cas_n
            sdram_wire_cke                                  : out   std_logic;                                        -- cke
            sdram_wire_cs_n                                 : out   std_logic;                                        -- cs_n
            sdram_wire_dq                                   : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
            sdram_wire_dqm                                  : out   std_logic_vector(1 downto 0);                     -- dqm
            sdram_wire_ras_n                                : out   std_logic;                                        -- ras_n
            sdram_wire_we_n                                 : out   std_logic;                                        -- we_n
            sdram_clk_clk                                   : out   std_logic;                                        -- clk
            sram_0_external_interface_DQ                    : inout std_logic_vector(15 downto 0) := (others => 'X'); -- DQ
            sram_0_external_interface_ADDR                  : out   std_logic_vector(17 downto 0);                    -- ADDR
            sram_0_external_interface_LB_N                  : out   std_logic;                                        -- LB_N
            sram_0_external_interface_UB_N                  : out   std_logic;                                        -- UB_N
            sram_0_external_interface_CE_N                  : out   std_logic;                                        -- CE_N
            sram_0_external_interface_OE_N                  : out   std_logic;                                        -- OE_N
            sram_0_external_interface_WE_N                  : out   std_logic;                                        -- WE_N
            video_vga_controller_0_external_interface_CLK   : out   std_logic;                                        -- CLK
            video_vga_controller_0_external_interface_HS    : out   std_logic;                                        -- HS
            video_vga_controller_0_external_interface_VS    : out   std_logic;                                        -- VS
            video_vga_controller_0_external_interface_BLANK : out   std_logic;                                        -- BLANK
            video_vga_controller_0_external_interface_SYNC  : out   std_logic;                                        -- SYNC
            video_vga_controller_0_external_interface_R     : out   std_logic_vector(9 downto 0);                     -- R
            video_vga_controller_0_external_interface_G     : out   std_logic_vector(9 downto 0);                     -- G
            video_vga_controller_0_external_interface_B     : out   std_logic_vector(9 downto 0)                      -- B
        );
    end component VGA_GRAPHICS;
		SIGNAL DQM : STD_LOGIC_VECTOR(1 DOWNTO 0);
		SIGNAL BA : STD_LOGIC_VECTOR(1 DOWNTO 0);
	BEGIN
		DRAM_BA_0 <= BA(0);
		DRAM_BA_1 <= BA(1);
		DRAM_UDQM <= DQM(1);
		DRAM_LDQM <= DQM(0);
	--instantiate NIOS II syste entity generated by the Qsys tool
		NiosII: VGA_GRAPHICS PORT MAP(
				clk_clk => CLOCK_50,
				reset_reset_n => KEY(0),
				sdram_clk_clk => DRAM_CLK,
				sdram_wire_addr => DRAM_ADDR,
				sdram_wire_ba => BA,
				sdram_wire_cas_n => DRAM_CAS_N,
				sdram_wire_cke => DRAM_CKE,
				sdram_wire_cs_n => DRAM_CS_N,
				sdram_wire_dq => DRAM_DQ,
				sdram_wire_dqm => DQM,
				sdram_wire_ras_n => DRAM_RAS_N,
				sdram_wire_we_n => DRAM_WE_N,
				
				video_vga_controller_0_external_interface_CLK	=>	VGA_CLK,	
				video_vga_controller_0_external_interface_HS	=>	VGA_HS,	
				video_vga_controller_0_external_interface_VS	=>	VGA_VS,	
				video_vga_controller_0_external_interface_BLANK	=>	VGA_BLANK,	
				video_vga_controller_0_external_interface_SYNC	=>	VGA_SYNC,	
				video_vga_controller_0_external_interface_R	=>	VGA_R,	
				video_vga_controller_0_external_interface_G	=>	VGA_G,	
				video_vga_controller_0_external_interface_B	=>	VGA_B,
				
				sram_0_external_interface_DQ	=>	SRAM_DQ,
				sram_0_external_interface_ADDR	=>	SRAM_ADDR,
				sram_0_external_interface_LB_N	=>	SRAM_LB_N,
				sram_0_external_interface_UB_N	=>	SRAM_UB_N,			
				sram_0_external_interface_CE_N	=>	SRAM_CE_N,
				sram_0_external_interface_OE_N	=>	SRAM_OE_N,
				sram_0_external_interface_WE_N	=>	SRAM_WE_N
			);
	END STRUCTURE;
	
	
